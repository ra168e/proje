asd
vehey
vehey_2