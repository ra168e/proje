asd
vehey
Vehey