asd
vehey